//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module parallel_to_serial
# (
    parameter width = 8
)
(
    input                      clk,
    input                      rst,

    input                      parallel_valid,
    input        [width - 1:0] parallel_data,

    output                     busy,
    output logic               serial_valid,
    output logic               serial_data
);
    // Task:
    // Implement a module that converts multi-bit parallel value to the single-bit serial data.
    //
    // The module should accept 'width' bit input parallel data when 'parallel_valid' input is asserted.
    // At the same clock cycle as 'parallel_valid' is asserted, the module should output
    // the least significant bit of the input data. In the following clock cycles the module
    // should output all the remaining bits of the parallel_data.
    // Together with providing correct 'serial_data' value, module should also assert the 'serial_valid' output.
    //
    // Note:
    // Check the waveform diagram in the README for better understanding.

    logic [width - 1:0] parallel_buffer;
    logic [$clog2(width):0] serial_counter;

    always_comb
    begin
        if(parallel_valid)
        begin
            serial_valid <= '1;
            serial_data <= parallel_data[0];
        end
        else if(serial_counter != 0)
        begin
            serial_valid <= '1;
            // busy = 1'b1;
            serial_data <= parallel_data[width-serial_counter];
        end
        else
        begin
            serial_valid <= '0;
            // busy = 1'b0;
        end

    end

    assign busy = serial_counter != 0 ? 1'b1 : 1'b0;

    always_ff @ (posedge clk)
    begin
        if(rst)
        begin
            parallel_buffer <= '0;
            serial_counter <= '0;
        end
        else if(parallel_valid)
        begin
            parallel_buffer <= parallel_data;
            serial_counter <= width-1;
        end
        else if(serial_counter > 0)
        begin
            serial_counter <= serial_counter - 1'b1;
        end
    end


endmodule
